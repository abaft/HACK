module mojo_top(
    // 50MHz clock input
    input clk,
    // Input from reset button (active low)
    input rst_n,
    // cclk input from AVR, high when AVR is ready
    input cclk,
    // Outputs to the 8 onboard LEDs
    output[7:0]led,
    // AVR SPI connections
    output spi_miso,
    input spi_ss,
    input spi_mosi,
    input spi_sck,
    // AVR ADC channel select
    output [3:0] spi_channel,
    // Serial connections
    input avr_tx, // AVR Tx => FPGA Rx
    output avr_rx, // AVR Rx => FPGA Tx
    input avr_rx_busy, // AVR Rx buffer full
    input [3:0] sw1,
	 input [3:0] sw2,
	 input [5:0] ctrl
	 );

wire rst = ~rst_n; // make reset active high

reg [7:0] LEDCTRL;

// these signals should be high-z when not used
assign spi_miso = 1'bz;
assign avr_rx = 1'bz;
assign spi_channel = 4'bzzzz;

//assign led = LEDCTRL;

reg [15:0] a = 16'b1101010001001110;
reg [15:0] b = 16'b0100101101101101;
reg c;

ALU(.x(sw1), .y(sw2), .control(ctrl), .out(led[3:0]), .zr(led[4]), .ng(led[5]));

endmodule